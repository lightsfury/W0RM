`timescale 1ns/100ps

module W0RM_Core_Branch #(
  parameter SINGLE_CYCLE = 0
)(
  input wire      clk
);

endmodule