`timescale 1ns/100ps

module W0RM_ALU_AddSub #(
  parameter SINGLE_CYCLE  = 0,
  parameter DATA_WIDTH    = 8
)(
  input wire                    clk,
  
  input wire                    data_valid,
  input wire  [3:0]             opcode,
  
  input wire  [DATA_WIDTH-1:0]  data_a,
                                data_b,
  
  output wire [DATA_WIDTH-1:0]  result,
  output wire                   result_valid,
  output wire [3:0]             result_flags
);
  localparam MSB            = DATA_WIDTH - 1;
  
  localparam ALU_OPCODE_ADD = 4'h8;
  localparam ALU_OPCODE_SUB = 4'h9;
  
  localparam ALU_FLAG_ZERO  = 4'h0;
  localparam ALU_FLAG_NEG   = 4'h1;
  localparam ALU_FLAG_OVER  = 4'h2;
  localparam ALU_FLAG_CARRY = 4'h3;
  
  reg   [DATA_WIDTH-1:0]  result_r = 0,
                          data_a_r = 0,
                          data_b_r = 0;
  reg                     flag_carry_r = 0,
                          flag_carry_i = 0,
                          result_valid_r = 0;
  reg   [DATA_WIDTH-1:0]  result_i = 0;
  
  assign result_flags[ALU_FLAG_ZERO]  = result_r == 0;
  assign result_flags[ALU_FLAG_NEG]   = result_r[MSB];
  assign result_flags[ALU_FLAG_OVER]  = ((~result_r[MSB]) && data_a_r[MSB] && data_b_r[MSB]) ||
                                        (result_r[MSB] && (~data_a_r[MSB]) && (~data_b_r[MSB]));
  assign result_flags[ALU_FLAG_CARRY] = flag_carry_r; // Carry generated by IP core
  
  assign result = result_r;
  assign result_valid = result_valid_r;
  
  always @(opcode, data_a, data_b)
  begin
    case (opcode)
      ALU_OPCODE_ADD:
        {flag_carry_i, result_i}  = (data_a + data_b);
      
      ALU_OPCODE_SUB:
        {flag_carry_i, result_i}  = (data_a + ~data_b) + 1;
      
      default:
      begin
        result_i      = {DATA_WIDTH{1'b0}};
        flag_carry_i  = 0;
      end
    endcase
  end
  
  generate
    if (SINGLE_CYCLE)
    begin
      
      always @(result_i, data_valid, data_a, data_b, flag_carry_i)
      begin
        result_r        = result_i;
        result_valid_r  = data_valid;
        data_a_r        = data_a;
        data_b_r        = data_b;
        flag_carry_r    = flag_carry_i;
      end
    end
    else
    begin
      always @(posedge clk)
      begin
        result_valid_r  <= data_valid;
        
        if (data_valid)
        begin
          data_a_r      <= data_a;
          data_b_r      <= data_b;
          
          result_r      <= result_i;
          flag_carry_r  <= flag_carry_i;
        end
      end
    end
  endgenerate
endmodule
