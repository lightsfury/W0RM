`timescale 1ns/100ps

module W0RM_Core_IFetch #(
  parameter SINGLE_CYCLE = 0
)(
  input wire      clk
);

endmodule