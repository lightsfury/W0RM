`timescale 1ns/100ps

module Visual_tests_tb(
  output wire done,
              error
);
  W0RM_Static_Timer_tb timer_tb();
  W0RM_Example_Design_tb();
  //Static_Timer_tb timer_tb;

endmodule
